module CSkA();
